// ------------------------------------------------------
//-------------------- тестовый набор  ------------------
// ------------------------------------------------------
parameter int ID_tag = 0;
parameter int Max_Burst_Len = 16;
parameter int RW_Delay_Value = 4;
parameter int Base_Address = 400;
parameter int Memory_Size = 100;
parameter int MIG_Port_Size = 128;
parameter int IO_Fifo_Depth = 32;
